module hello

pub fn hello() string {
	return 'Hello, '
}
