module hello

fn test_hello() {
	assert hello() == 'Hello, '
}
